`timescale 1ns/1ps

module mailbox_example;

endmodule

